import_C( "cygwin_tecs.h" );

signature sSample {
  ER  sayHello( [in]int32_t times );
  ER  howAreYou( [out, string(len)]char_t *buf, [in]int32_t len );
};

celltype tSample {
  entry sSample eEnt;
};

celltype tSimple {
  call sSample cCall;
  entry sTaskBody eBody;
};

cell tSample Sample {
};

cell tSimple Simple {
  cCall = Sample.eEnt;
};

cell tTask Task {
  cBody = Simple.eBody;
  priority = 11;
  stackSize = 1024;
  taskAttribute = C_EXP( "TA_AcT" );
};