import_C("ev3api_motor.h");
signature sMotor{
	ER_UINT getType(void);
	int32_t getCounts(void);
	int getPower(void);
	ER resetCounts(void);
	ER setPower([in]int power);
	ER stop([in] bool_t brake); 
	ER rotate([in] int degrees, [in] uint32_t speed_abs, [in]bool_t blocking);
	// ER ev3_motor_steer(motor_port_t left_motor, motor_port_t right_motor, int power, int turn_ratio);
	void initializePort([in]int32_t type);
};

celltype tMotor{
	entry sMotor eMotor;
	attr{
		int32_t port;
	};
};
